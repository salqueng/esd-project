module Logic_out (High, Low, Z);
	output High, Low, Z;
	
	assign High = 1'b1;
	assign Low  = 1'b0;
	assign Z    = 1'bz;
endmodule
